��G.      �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�	estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �_sklearn_version��1.2.2�ub�n_estimators�K
�estimator_params�(hhhhhhhhhht��base_estimator��
deprecated��	bootstrap���	oob_score���n_jobs�NhK �verbose�K �
warm_start��hN�max_samples�NhhhKhKhKhG        h�sqrt�hNhG        hG        �feature_names_in_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h+�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�objawy��wiek��choroby_wsp��wzrost��leki�et�b�n_features_in_�K�
n_outputs_�K�classes_�h*h-K ��h/��R�(KK��h4�i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�
n_classes_�K�
estimator_�h	�estimators_�]�(h)��}�(hhhhhKhKhKhG        hh&hNhJ�
hG        hNhG        hAKhBKhCh*h-K ��h/��R�(KK��h4�f8�����R�(KhKNNNJ����J����K t�b�C              �?�t�bhOh(�scalar���hJC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���Kh*h-K ��h/��R�(KK��hJ�C       �t�bK��R�}�(hK�
node_count�K�nodes�h*h-K ��h/��R�(KK��h4�V56�����R�(Kh8N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(h{h4�i8�����R�(KhKNNNJ����J����K t�bK ��h|h�K��h}h�K��h~h[K��hh[K ��h�h�K(��h�h[K0��uK8KKt�b�B�                             �?r�qG�?             H@                           �?      �?	             0@������������������������       �                     @                            �?�<ݚ�?             "@������������������������       �                     @������������������������       ����Q��?             @       
                   �g@     ��?             @@       	                    @�t����?             1@������������������������       �                     $@������������������������       �����X�?             @                           @�r����?             .@������������������������       �z�G�z�?             $@������������������������       �                     @�t�b�values�h*h-K ��h/��R�(KKKK��h[�C�      ?@      1@      ,@       @      @              @       @      @              @       @      1@      .@      .@       @      $@              @       @       @      *@       @       @              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh&hNhJ/��hG        hNhG        hAKhBKhCh*h-K ��h/��R�(KK��h[�C              �?�t�bhOh`hJC       ���R�hdKhehhKh*h-K ��h/��R�(KK��hJ�C       �t�bK��R�}�(hKhrKhsh*h-K ��h/��R�(KK��hz�Bh                            �g@r�q��?!             H@                          �E@f���M�?             ?@                          �e@b�2�tk�?             2@������������������������       �      �?              @������������������������       �z�G�z�?             $@������������������������       �                     *@       
                     @�t����?             1@       	                    �?      �?              @������������������������       �؇���X�?             @������������������������       �                     �?������������������������       �                     "@�t�bh�h*h-K ��h/��R�(KKKK��h[�C�      6@      :@      4@      &@      @      &@      @      @       @       @      *@               @      .@       @      @      �?      @      �?                      "@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh&hNhJu�7hG        hNhG        hAKhBKhCh*h-K ��h/��R�(KK��h[�C              �?�t�bhOh`hJC       ���R�hdKhehhKh*h-K ��h/��R�(KK��hJ�C       �t�bK��R�}�(hKhrKhsh*h-K ��h/��R�(KK��hz�Bh                            @K@     ��?             H@                           �?"pc�
�?            �@@������������������������       �                     @                          �T@�θ�?             :@������������������������       �                     �?������������������������       �z�G�z�?             9@       
                   Ph@���Q��?             .@       	                     @"pc�
�?             &@������������������������       �                     @������������������������       �      �?             @������������������������       �                     @�t�bh�h*h-K ��h/��R�(KKKK��h[�C�      .@     �@@      @      ;@              @      @      4@      �?              @      4@      "@      @      "@       @      @               @       @              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh&hNhJ��!XhG        hNhG        hAKhBKhCh*h-K ��h/��R�(KK��h[�C              �?�t�bhOh`hJC       ���R�hdKhehhKh*h-K ��h/��R�(KK��hJ�C       �t�bK��R�}�(hKhrK	hsh*h-K ��h/��R�(KK	��hz�B�                              �?�q���?             H@                          �g@      �?             0@������������������������       �                     ,@������������������������       �                      @                           @     ��?             @@                          �f@
j*D>�?             :@������������������������       �X�Cc�?	             ,@������������������������       �r�q��?             (@������������������������       �                     @�t�bh�h*h-K ��h/��R�(KK	KK��h[�C�      9@      7@      ,@       @      ,@                       @      &@      5@      &@      .@      "@      @       @      $@              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh&hNhJC�NhG        hNhG        hAKhBKhCh*h-K ��h/��R�(KK��h[�C              �?�t�bhOh`hJC       ���R�hdKhehhKh*h-K ��h/��R�(KK��hJ�C       �t�bK��R�}�(hKhrKhsh*h-K ��h/��R�(KK��hz�Bh                             �?�q���?#             H@                          �E@�����?             3@                           @և���X�?
             ,@������������������������       �                     @������������������������       ��eP*L��?             &@������������������������       �                     @       
                     @�f7�z�?             =@       	                   �C@�q�����?             9@������������������������       �      �?	             (@������������������������       ��	j*D�?             *@������������������������       �                     @�t�bh�h*h-K ��h/��R�(KKKK��h[�C�      9@      7@      *@      @       @      @      @              @      @      @              (@      1@      (@      *@      @      "@      "@      @              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh&hNhJ�R�[hG        hNhG        hAKhBKhCh*h-K ��h/��R�(KK��h[�C              �?�t�bhOh`hJC       ���R�hdKhehhKh*h-K ��h/��R�(KK��hJ�C       �t�bK��R�}�(hKhrKhsh*h-K ��h/��R�(KK��hz�Bh                            �E@     ��?             H@                          �e@�q�q�?             8@                           @���Q��?             @������������������������       �                      @������������������������       ��q�q�?             @                           @���y4F�?             3@������������������������       �                     @������������������������       �����X�?
             ,@	       
                   0h@r�q��?             8@������������������������       �        	             4@������������������������       �                     @�t�bh�h*h-K ��h/��R�(KKKK��h[�C�      ;@      5@      @      1@      @       @       @              �?       @      @      .@              @      @      $@      4@      @      4@                      @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh&hNhJ�v}hG        hNhG        hAKhBKhCh*h-K ��h/��R�(KK��h[�C              �?�t�bhOh`hJC       ���R�hdKhehhKh*h-K ��h/��R�(KK��hJ�C       �t�bK��R�}�(hKhrKhsh*h-K ��h/��R�(KK��hz�B�                            �E@      �?             H@                          �0@4�2%ޑ�?            �A@                          `f@      �?              @������������������������       �                     @������������������������       ����Q��?             @                           6@�>����?             ;@������������������������       �r�q��?             @������������������������       ����N8�?             5@	                          �Q@�θ�?	             *@
                          �g@r�q��?             (@������������������������       �                      @������������������������       �      �?             @������������������������       �                     �?�t�bh�h*h-K ��h/��R�(KKKK��h[�C�      2@      >@       @      ;@      @       @      @              @       @       @      9@      �?      @      �?      4@      $@      @      $@       @       @               @       @              �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh&hNhJg}�XhG        hNhG        hAKhBKhCh*h-K ��h/��R�(KK��h[�C              �?�t�bhOh`hJC       ���R�hdKhehhKh*h-K ��h/��R�(KK��hJ�C       �t�bK��R�}�(hKhrKhsh*h-K ��h/��R�(KK��hz�B�                            �g@�q�q�?             H@                            @�<ݚ�?             B@                          �e@z�G�z�?            �A@������������������������       �ףp=
�?             4@������������������������       ��q�q�?
             .@������������������������       �                     �?������������������������       �                     (@�t�bh�h*h-K ��h/��R�(KKKK��h[�Cp      <@      4@      <@       @      <@      @      2@       @      $@      @              �?              (@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh&hNhJ	�tlhG        hNhG        hAKhBKhCh*h-K ��h/��R�(KK��h[�C              �?�t�bhOh`hJC       ���R�hdKhehhKh*h-K ��h/��R�(KK��hJ�C       �t�bK��R�}�(hKhrK	hsh*h-K ��h/��R�(KK	��hz�B�                              �?      �?             H@������������������������       �                     &@                          pg@^H���+�?            �B@                            @      �?             0@������������������������       ��q�q�?             .@������������������������       �                     �?                           7@؇���X�?             5@������������������������       ����Q��?             @������������������������       �      �?
             0@�t�bh�h*h-K ��h/��R�(KK	KK��h[�C�      8@      8@      &@              *@      8@      $@      @      $@      @              �?      @      2@       @      @      �?      .@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh&hNhJ�ޡhG        hNhG        hAKhBKhCh*h-K ��h/��R�(KK��h[�C              �?�t�bhOh`hJC       ���R�hdKhehhKh*h-K ��h/��R�(KK��hJ�C       �t�bK��R�}�(hKhrK	hsh*h-K ��h/��R�(KK	��hz�B�                              �?      �?             H@������������������������       �                     ,@                            @��.k���?             A@                          �0@�	j*D�?	             *@������������������������       ��q�q�?             @������������������������       �                     @                           @և���X�?             5@������������������������       �z�G�z�?             .@������������������������       �                     @�t�bh�h*h-K ��h/��R�(KK	KK��h[�C�      >@      2@      ,@              0@      2@      @      "@      @       @              @      (@      "@      (@      @              @�t�bubhhubehhub.